`timescale 1ns/1ns

module bothmult(input [5:0] inbus,
           input start, clk, rst,
           output [5:0] outbus,
           output ready);
        

  wire [1:0] decision_bits ;
  wire ldX, ldY, lde, ldA, shA, shX, clrA, clrX, clre,
      add, sub;
  wire [1:0] upload_selector;
  logic finished;
  controller cu(clk, rst, start, decision_bits,ldX, ldY, lde, ldA, shA, shX, clrA, clrX, clre,
      add, sub ,finished, upload_selector);
  dataPath dp(inbus, ldX, shX, clrX , ldY, ldA, shA, clrA, lde, clre, add, sub, clk, rst, upload_selector, outbus, decision_bits);
  assign ready = finished;
endmodule
