`timescale 1ns/1ns

module b1reg (input in, clr, load, clk, rst, output reg out);
  always@(posedge clk, posedge rst)begin
    if(rst)
      out = 1'b0;
    else
      if(clr)
        out = 1'b0;
      else
        if(load)
          out <= in;
  end
endmodule

